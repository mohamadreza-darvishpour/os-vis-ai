-------------------------------------------------------------------------------
--
-- Title       : TrafficLightController_tb
-- Design      : sys_dig_des
-- Author      : fardad
-- Company     : .
--
-------------------------------------------------------------------------------
--
-- File        : C:\Users\beta\Documents\0-parseh-ai-os-vis\z_digital_system\active_hdl\my_project_files\TrafficLightController_Workspace\sys_dig_des\src\TrafficLightController_tb.vhd
-- Generated   : Fri Dec 27 17:43:18 2024
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {TrafficLightController_tb} architecture {TrafficLightController_tb}}

library IEEE;
use IEEE.std_logic_1164.all;

entity TrafficLightController_tb is
	 port(
		 Y1 : out STD_LOGIC;
		 Y2 : out STD_LOGIC;
		 G1 : out STD_LOGIC;
		 G2 : out STD_LOGIC;
		 R1 : out STD_LOGIC;
		 R2 : out STD_LOGIC;
		 clk : in STD_LOGIC
	     );
end TrafficLightController_tb;

--}} End of automatically maintained section

architecture TrafficLightController_tb of TrafficLightController_tb is
begin

	 -- enter your statements here --

end TrafficLightController_tb;
